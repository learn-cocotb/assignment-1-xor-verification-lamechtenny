module exor_text(
                input wire a,b,
                output wire y);
exor
